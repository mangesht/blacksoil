if ($value$plusargs("TESTNAME=%s", testname)) begin
    $display("Running test %0s.", testname);
  startTest();
end 

