Lets keep somethings 