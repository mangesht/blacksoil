covergroup hdrTransitions;
coverpoint tempHdr {
    bins EthIpv4TcpTrans = (Eth =>Ipv4 =>Tcp);
    bins EthIpv6TcpTrans = (Eth =>Ipv6 =>Tcp);
    bins EthIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMpls1InnerIpv4Trans = (Eth =>Mpls1 =>InnerIpv4);
    bins EthMpls1InnerIpv6Trans = (Eth =>Mpls1 =>InnerIpv6);
    bins EthMpls1InnerEthTrans = (Eth =>Mpls1 =>InnerEth);
    bins EthMpls1Mpls2InnerIpv4Trans = (Eth =>Mpls1Mpls2 =>InnerIpv4);
    bins EthMpls1Mpls2InnerIpv6Trans = (Eth =>Mpls1Mpls2 =>InnerIpv6);
    bins EthMpls1Mpls2InnerEthTrans = (Eth =>Mpls1Mpls2 =>InnerEth);
    bins EthMpls1Mpls2Mpls3InnerIpv4Trans = (Eth =>Mpls1Mpls2Mpls3 =>InnerIpv4);
    bins EthMpls1Mpls2Mpls3InnerIpv6Trans = (Eth =>Mpls1Mpls2Mpls3 =>InnerIpv6);
    bins EthMpls1Mpls2Mpls3InnerEthTrans = (Eth =>Mpls1Mpls2Mpls3 =>InnerEth);
    bins EthL2SiaIpv4TcpTrans = (Eth =>L2Sia =>Ipv4 =>Tcp);
    bins EthL2SiaIpv6TcpTrans = (Eth =>L2Sia =>Ipv6 =>Tcp);
    bins EthL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthL2SiaMpls1InnerIpv4Trans = (Eth =>L2Sia =>Mpls1 =>InnerIpv4);
    bins EthL2SiaMpls1InnerIpv6Trans = (Eth =>L2Sia =>Mpls1 =>InnerIpv6);
    bins EthL2SiaMpls1InnerEthTrans = (Eth =>L2Sia =>Mpls1 =>InnerEth);
    bins EthL2SiaMpls1Mpls2InnerIpv4Trans = (Eth =>L2Sia =>Mpls1Mpls2 =>InnerIpv4);
    bins EthL2SiaMpls1Mpls2InnerIpv6Trans = (Eth =>L2Sia =>Mpls1Mpls2 =>InnerIpv6);
    bins EthL2SiaMpls1Mpls2InnerEthTrans = (Eth =>L2Sia =>Mpls1Mpls2 =>InnerEth);
    bins EthL2SiaMpls1Mpls2Mpls3InnerIpv4Trans = (Eth =>L2Sia =>Mpls1Mpls2Mpls3 =>InnerIpv4);
    bins EthL2SiaMpls1Mpls2Mpls3InnerIpv6Trans = (Eth =>L2Sia =>Mpls1Mpls2Mpls3 =>InnerIpv6);
    bins EthL2SiaMpls1Mpls2Mpls3InnerEthTrans = (Eth =>L2Sia =>Mpls1Mpls2Mpls3 =>InnerEth);
    bins EthTag1qIpv4TcpTrans = (Eth =>Tag1q =>Ipv4 =>Tcp);
    bins EthTag1qIpv6TcpTrans = (Eth =>Tag1q =>Ipv6 =>Tcp);
    bins EthTag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>Tag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthTag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>Tag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthTag1qL2SiaIpv4TcpTrans = (Eth =>Tag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthTag1qL2SiaIpv6TcpTrans = (Eth =>Tag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthTag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>Tag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthTag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>Tag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthTag1qTag1qIpv4TcpTrans = (Eth =>Tag1qTag1q =>Ipv4 =>Tcp);
    bins EthTag1qTag1qIpv6TcpTrans = (Eth =>Tag1qTag1q =>Ipv6 =>Tcp);
    bins EthTag1qTag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>Tag1qTag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthTag1qTag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>Tag1qTag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthTag1qTag1qL2SiaIpv4TcpTrans = (Eth =>Tag1qTag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthTag1qTag1qL2SiaIpv6TcpTrans = (Eth =>Tag1qTag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthTag1qTag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>Tag1qTag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthTag1qTag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>Tag1qTag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthStagIpv4TcpTrans = (Eth =>Stag =>Ipv4 =>Tcp);
    bins EthStagIpv6TcpTrans = (Eth =>Stag =>Ipv6 =>Tcp);
    bins EthStagIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>Stag =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthStagIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>Stag =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthStagL2SiaIpv4TcpTrans = (Eth =>Stag =>L2Sia =>Ipv4 =>Tcp);
    bins EthStagL2SiaIpv6TcpTrans = (Eth =>Stag =>L2Sia =>Ipv6 =>Tcp);
    bins EthStagL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>Stag =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthStagL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>Stag =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthStagTag1qIpv4TcpTrans = (Eth =>StagTag1q =>Ipv4 =>Tcp);
    bins EthStagTag1qIpv6TcpTrans = (Eth =>StagTag1q =>Ipv6 =>Tcp);
    bins EthStagTag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>StagTag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthStagTag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>StagTag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthStagTag1qL2SiaIpv4TcpTrans = (Eth =>StagTag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthStagTag1qL2SiaIpv6TcpTrans = (Eth =>StagTag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthStagTag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>StagTag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthStagTag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>StagTag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthVnTagTag1qIpv4TcpTrans = (Eth =>VnTag =>Tag1q =>Ipv4 =>Tcp);
    bins EthVnTagTag1qIpv6TcpTrans = (Eth =>VnTag =>Tag1q =>Ipv6 =>Tcp);
    bins EthVnTagTag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>VnTag =>Tag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthVnTagTag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>VnTag =>Tag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthVnTagTag1qL2SiaIpv4TcpTrans = (Eth =>VnTag =>Tag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthVnTagTag1qL2SiaIpv6TcpTrans = (Eth =>VnTag =>Tag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthVnTagTag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>VnTag =>Tag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthVnTagTag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>VnTag =>Tag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthVnTagTag1qL2CmdIpv4TcpTrans = (Eth =>VnTag =>Tag1q =>L2Cmd =>Ipv4 =>Tcp);
    bins EthVnTagTag1qL2CmdIpv6TcpTrans = (Eth =>VnTag =>Tag1q =>L2Cmd =>Ipv6 =>Tcp);
    bins EthVnTagTag1qL2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>VnTag =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthVnTagTag1qL2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>VnTag =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthVnTagTag1qL2CmdL2SiaIpv4TcpTrans = (Eth =>VnTag =>Tag1q =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthVnTagTag1qL2CmdL2SiaIpv6TcpTrans = (Eth =>VnTag =>Tag1q =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthVnTagTag1qL2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>VnTag =>Tag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthVnTagTag1qL2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>VnTag =>Tag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthVnTagTag1qTag1qIpv4TcpTrans = (Eth =>VnTag =>Tag1qTag1q =>Ipv4 =>Tcp);
    bins EthVnTagTag1qTag1qIpv6TcpTrans = (Eth =>VnTag =>Tag1qTag1q =>Ipv6 =>Tcp);
    bins EthVnTagTag1qTag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>VnTag =>Tag1qTag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthVnTagTag1qTag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>VnTag =>Tag1qTag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthVnTagTag1qTag1qL2SiaIpv4TcpTrans = (Eth =>VnTag =>Tag1qTag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthVnTagTag1qTag1qL2SiaIpv6TcpTrans = (Eth =>VnTag =>Tag1qTag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthVnTagTag1qTag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>VnTag =>Tag1qTag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthVnTagTag1qTag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>VnTag =>Tag1qTag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthVnTagTag1qTag1qL2CmdIpv4TcpTrans = (Eth =>VnTag =>Tag1qTag1q =>L2Cmd =>Ipv4 =>Tcp);
    bins EthVnTagTag1qTag1qL2CmdIpv6TcpTrans = (Eth =>VnTag =>Tag1qTag1q =>L2Cmd =>Ipv6 =>Tcp);
    bins EthVnTagTag1qTag1qL2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>VnTag =>Tag1qTag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthVnTagTag1qTag1qL2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>VnTag =>Tag1qTag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthVnTagTag1qTag1qL2CmdL2SiaIpv4TcpTrans = (Eth =>VnTag =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthVnTagTag1qTag1qL2CmdL2SiaIpv6TcpTrans = (Eth =>VnTag =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthVnTagTag1qTag1qL2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>VnTag =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthVnTagTag1qTag1qL2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>VnTag =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthVnTagStagTag1qIpv4TcpTrans = (Eth =>VnTag =>StagTag1q =>Ipv4 =>Tcp);
    bins EthVnTagStagTag1qIpv6TcpTrans = (Eth =>VnTag =>StagTag1q =>Ipv6 =>Tcp);
    bins EthVnTagStagTag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>VnTag =>StagTag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthVnTagStagTag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>VnTag =>StagTag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthVnTagStagTag1qL2SiaIpv4TcpTrans = (Eth =>VnTag =>StagTag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthVnTagStagTag1qL2SiaIpv6TcpTrans = (Eth =>VnTag =>StagTag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthVnTagStagTag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>VnTag =>StagTag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthVnTagStagTag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>VnTag =>StagTag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthVnTagStagTag1qL2CmdIpv4TcpTrans = (Eth =>VnTag =>StagTag1q =>L2Cmd =>Ipv4 =>Tcp);
    bins EthVnTagStagTag1qL2CmdIpv6TcpTrans = (Eth =>VnTag =>StagTag1q =>L2Cmd =>Ipv6 =>Tcp);
    bins EthVnTagStagTag1qL2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>VnTag =>StagTag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthVnTagStagTag1qL2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>VnTag =>StagTag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthVnTagStagTag1qL2CmdL2SiaIpv4TcpTrans = (Eth =>VnTag =>StagTag1q =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthVnTagStagTag1qL2CmdL2SiaIpv6TcpTrans = (Eth =>VnTag =>StagTag1q =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthVnTagStagTag1qL2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>VnTag =>StagTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthVnTagStagTag1qL2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>VnTag =>StagTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthSilTag1qIpv4TcpTrans = (Eth =>Sil =>Tag1q =>Ipv4 =>Tcp);
    bins EthSilTag1qIpv6TcpTrans = (Eth =>Sil =>Tag1q =>Ipv6 =>Tcp);
    bins EthSilTag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>Sil =>Tag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthSilTag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>Sil =>Tag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthSilTag1qL2SiaIpv4TcpTrans = (Eth =>Sil =>Tag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthSilTag1qL2SiaIpv6TcpTrans = (Eth =>Sil =>Tag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthSilTag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>Sil =>Tag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthSilTag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>Sil =>Tag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthSilTag1qL2CmdIpv4TcpTrans = (Eth =>Sil =>Tag1q =>L2Cmd =>Ipv4 =>Tcp);
    bins EthSilTag1qL2CmdIpv6TcpTrans = (Eth =>Sil =>Tag1q =>L2Cmd =>Ipv6 =>Tcp);
    bins EthSilTag1qL2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>Sil =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthSilTag1qL2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>Sil =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthSilTag1qL2CmdL2SiaIpv4TcpTrans = (Eth =>Sil =>Tag1q =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthSilTag1qL2CmdL2SiaIpv6TcpTrans = (Eth =>Sil =>Tag1q =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthSilTag1qL2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>Sil =>Tag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthSilTag1qL2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>Sil =>Tag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthSilTag1qTag1qIpv4TcpTrans = (Eth =>Sil =>Tag1qTag1q =>Ipv4 =>Tcp);
    bins EthSilTag1qTag1qIpv6TcpTrans = (Eth =>Sil =>Tag1qTag1q =>Ipv6 =>Tcp);
    bins EthSilTag1qTag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>Sil =>Tag1qTag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthSilTag1qTag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>Sil =>Tag1qTag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthSilTag1qTag1qL2SiaIpv4TcpTrans = (Eth =>Sil =>Tag1qTag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthSilTag1qTag1qL2SiaIpv6TcpTrans = (Eth =>Sil =>Tag1qTag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthSilTag1qTag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>Sil =>Tag1qTag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthSilTag1qTag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>Sil =>Tag1qTag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthSilTag1qTag1qL2CmdIpv4TcpTrans = (Eth =>Sil =>Tag1qTag1q =>L2Cmd =>Ipv4 =>Tcp);
    bins EthSilTag1qTag1qL2CmdIpv6TcpTrans = (Eth =>Sil =>Tag1qTag1q =>L2Cmd =>Ipv6 =>Tcp);
    bins EthSilTag1qTag1qL2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>Sil =>Tag1qTag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthSilTag1qTag1qL2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>Sil =>Tag1qTag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthSilTag1qTag1qL2CmdL2SiaIpv4TcpTrans = (Eth =>Sil =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthSilTag1qTag1qL2CmdL2SiaIpv6TcpTrans = (Eth =>Sil =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthSilTag1qTag1qL2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>Sil =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthSilTag1qTag1qL2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>Sil =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthSilVnTagTag1qIpv4TcpTrans = (Eth =>Sil =>VnTag =>Tag1q =>Ipv4 =>Tcp);
    bins EthSilVnTagTag1qIpv6TcpTrans = (Eth =>Sil =>VnTag =>Tag1q =>Ipv6 =>Tcp);
    bins EthSilVnTagTag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>Sil =>VnTag =>Tag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthSilVnTagTag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>Sil =>VnTag =>Tag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthSilVnTagTag1qL2SiaIpv4TcpTrans = (Eth =>Sil =>VnTag =>Tag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthSilVnTagTag1qL2SiaIpv6TcpTrans = (Eth =>Sil =>VnTag =>Tag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthSilVnTagTag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>Sil =>VnTag =>Tag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthSilVnTagTag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>Sil =>VnTag =>Tag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthSilVnTagTag1qL2CmdIpv4TcpTrans = (Eth =>Sil =>VnTag =>Tag1q =>L2Cmd =>Ipv4 =>Tcp);
    bins EthSilVnTagTag1qL2CmdIpv6TcpTrans = (Eth =>Sil =>VnTag =>Tag1q =>L2Cmd =>Ipv6 =>Tcp);
    bins EthSilVnTagTag1qL2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>Sil =>VnTag =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthSilVnTagTag1qL2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>Sil =>VnTag =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthSilVnTagTag1qL2CmdL2SiaIpv4TcpTrans = (Eth =>Sil =>VnTag =>Tag1q =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthSilVnTagTag1qL2CmdL2SiaIpv6TcpTrans = (Eth =>Sil =>VnTag =>Tag1q =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthSilVnTagTag1qL2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>Sil =>VnTag =>Tag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthSilVnTagTag1qL2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>Sil =>VnTag =>Tag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthSilVnTagTag1qTag1qIpv4TcpTrans = (Eth =>Sil =>VnTag =>Tag1qTag1q =>Ipv4 =>Tcp);
    bins EthSilVnTagTag1qTag1qIpv6TcpTrans = (Eth =>Sil =>VnTag =>Tag1qTag1q =>Ipv6 =>Tcp);
    bins EthSilVnTagTag1qTag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>Sil =>VnTag =>Tag1qTag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthSilVnTagTag1qTag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>Sil =>VnTag =>Tag1qTag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthSilVnTagTag1qTag1qL2SiaIpv4TcpTrans = (Eth =>Sil =>VnTag =>Tag1qTag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthSilVnTagTag1qTag1qL2SiaIpv6TcpTrans = (Eth =>Sil =>VnTag =>Tag1qTag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthSilVnTagTag1qTag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>Sil =>VnTag =>Tag1qTag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthSilVnTagTag1qTag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>Sil =>VnTag =>Tag1qTag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthSilVnTagTag1qTag1qL2CmdIpv4TcpTrans = (Eth =>Sil =>VnTag =>Tag1qTag1q =>L2Cmd =>Ipv4 =>Tcp);
    bins EthSilVnTagTag1qTag1qL2CmdIpv6TcpTrans = (Eth =>Sil =>VnTag =>Tag1qTag1q =>L2Cmd =>Ipv6 =>Tcp);
    bins EthSilVnTagTag1qTag1qL2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>Sil =>VnTag =>Tag1qTag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthSilVnTagTag1qTag1qL2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>Sil =>VnTag =>Tag1qTag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthSilVnTagTag1qTag1qL2CmdL2SiaIpv4TcpTrans = (Eth =>Sil =>VnTag =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthSilVnTagTag1qTag1qL2CmdL2SiaIpv6TcpTrans = (Eth =>Sil =>VnTag =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthSilVnTagTag1qTag1qL2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>Sil =>VnTag =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthSilVnTagTag1qTag1qL2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>Sil =>VnTag =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8Ipv4TcpTrans = (Eth =>MacSec8 =>Ipv4 =>Tcp);
    bins EthMacSec8Ipv6TcpTrans = (Eth =>MacSec8 =>Ipv6 =>Tcp);
    bins EthMacSec8Ipv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8Ipv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8Mpls1InnerIpv4Trans = (Eth =>MacSec8 =>Mpls1 =>InnerIpv4);
    bins EthMacSec8Mpls1InnerIpv6Trans = (Eth =>MacSec8 =>Mpls1 =>InnerIpv6);
    bins EthMacSec8Mpls1InnerEthTrans = (Eth =>MacSec8 =>Mpls1 =>InnerEth);
    bins EthMacSec8Mpls1Mpls2InnerIpv4Trans = (Eth =>MacSec8 =>Mpls1Mpls2 =>InnerIpv4);
    bins EthMacSec8Mpls1Mpls2InnerIpv6Trans = (Eth =>MacSec8 =>Mpls1Mpls2 =>InnerIpv6);
    bins EthMacSec8Mpls1Mpls2InnerEthTrans = (Eth =>MacSec8 =>Mpls1Mpls2 =>InnerEth);
    bins EthMacSec8Mpls1Mpls2Mpls3InnerIpv4Trans = (Eth =>MacSec8 =>Mpls1Mpls2Mpls3 =>InnerIpv4);
    bins EthMacSec8Mpls1Mpls2Mpls3InnerIpv6Trans = (Eth =>MacSec8 =>Mpls1Mpls2Mpls3 =>InnerIpv6);
    bins EthMacSec8Mpls1Mpls2Mpls3InnerEthTrans = (Eth =>MacSec8 =>Mpls1Mpls2Mpls3 =>InnerEth);
    bins EthMacSec8L2SiaIpv4TcpTrans = (Eth =>MacSec8 =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec8L2SiaIpv6TcpTrans = (Eth =>MacSec8 =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec8L2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8L2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8L2SiaMpls1InnerIpv4Trans = (Eth =>MacSec8 =>L2Sia =>Mpls1 =>InnerIpv4);
    bins EthMacSec8L2SiaMpls1InnerIpv6Trans = (Eth =>MacSec8 =>L2Sia =>Mpls1 =>InnerIpv6);
    bins EthMacSec8L2SiaMpls1InnerEthTrans = (Eth =>MacSec8 =>L2Sia =>Mpls1 =>InnerEth);
    bins EthMacSec8L2SiaMpls1Mpls2InnerIpv4Trans = (Eth =>MacSec8 =>L2Sia =>Mpls1Mpls2 =>InnerIpv4);
    bins EthMacSec8L2SiaMpls1Mpls2InnerIpv6Trans = (Eth =>MacSec8 =>L2Sia =>Mpls1Mpls2 =>InnerIpv6);
    bins EthMacSec8L2SiaMpls1Mpls2InnerEthTrans = (Eth =>MacSec8 =>L2Sia =>Mpls1Mpls2 =>InnerEth);
    bins EthMacSec8L2SiaMpls1Mpls2Mpls3InnerIpv4Trans = (Eth =>MacSec8 =>L2Sia =>Mpls1Mpls2Mpls3 =>InnerIpv4);
    bins EthMacSec8L2SiaMpls1Mpls2Mpls3InnerIpv6Trans = (Eth =>MacSec8 =>L2Sia =>Mpls1Mpls2Mpls3 =>InnerIpv6);
    bins EthMacSec8L2SiaMpls1Mpls2Mpls3InnerEthTrans = (Eth =>MacSec8 =>L2Sia =>Mpls1Mpls2Mpls3 =>InnerEth);
    bins EthMacSec8L2CmdIpv4TcpTrans = (Eth =>MacSec8 =>L2Cmd =>Ipv4 =>Tcp);
    bins EthMacSec8L2CmdIpv6TcpTrans = (Eth =>MacSec8 =>L2Cmd =>Ipv6 =>Tcp);
    bins EthMacSec8L2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8L2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8L2CmdMpls1InnerIpv4Trans = (Eth =>MacSec8 =>L2Cmd =>Mpls1 =>InnerIpv4);
    bins EthMacSec8L2CmdMpls1InnerIpv6Trans = (Eth =>MacSec8 =>L2Cmd =>Mpls1 =>InnerIpv6);
    bins EthMacSec8L2CmdMpls1InnerEthTrans = (Eth =>MacSec8 =>L2Cmd =>Mpls1 =>InnerEth);
    bins EthMacSec8L2CmdMpls1Mpls2InnerIpv4Trans = (Eth =>MacSec8 =>L2Cmd =>Mpls1Mpls2 =>InnerIpv4);
    bins EthMacSec8L2CmdMpls1Mpls2InnerIpv6Trans = (Eth =>MacSec8 =>L2Cmd =>Mpls1Mpls2 =>InnerIpv6);
    bins EthMacSec8L2CmdMpls1Mpls2InnerEthTrans = (Eth =>MacSec8 =>L2Cmd =>Mpls1Mpls2 =>InnerEth);
    bins EthMacSec8L2CmdMpls1Mpls2Mpls3InnerIpv4Trans = (Eth =>MacSec8 =>L2Cmd =>Mpls1Mpls2Mpls3 =>InnerIpv4);
    bins EthMacSec8L2CmdMpls1Mpls2Mpls3InnerIpv6Trans = (Eth =>MacSec8 =>L2Cmd =>Mpls1Mpls2Mpls3 =>InnerIpv6);
    bins EthMacSec8L2CmdMpls1Mpls2Mpls3InnerEthTrans = (Eth =>MacSec8 =>L2Cmd =>Mpls1Mpls2Mpls3 =>InnerEth);
    bins EthMacSec8L2CmdL2SiaIpv4TcpTrans = (Eth =>MacSec8 =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec8L2CmdL2SiaIpv6TcpTrans = (Eth =>MacSec8 =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec8L2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8L2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8L2CmdL2SiaMpls1InnerIpv4Trans = (Eth =>MacSec8 =>L2Cmd =>L2Sia =>Mpls1 =>InnerIpv4);
    bins EthMacSec8L2CmdL2SiaMpls1InnerIpv6Trans = (Eth =>MacSec8 =>L2Cmd =>L2Sia =>Mpls1 =>InnerIpv6);
    bins EthMacSec8L2CmdL2SiaMpls1InnerEthTrans = (Eth =>MacSec8 =>L2Cmd =>L2Sia =>Mpls1 =>InnerEth);
    bins EthMacSec8L2CmdL2SiaMpls1Mpls2InnerIpv4Trans = (Eth =>MacSec8 =>L2Cmd =>L2Sia =>Mpls1Mpls2 =>InnerIpv4);
    bins EthMacSec8L2CmdL2SiaMpls1Mpls2InnerIpv6Trans = (Eth =>MacSec8 =>L2Cmd =>L2Sia =>Mpls1Mpls2 =>InnerIpv6);
    bins EthMacSec8L2CmdL2SiaMpls1Mpls2InnerEthTrans = (Eth =>MacSec8 =>L2Cmd =>L2Sia =>Mpls1Mpls2 =>InnerEth);
    bins EthMacSec8L2CmdL2SiaMpls1Mpls2Mpls3InnerIpv4Trans = (Eth =>MacSec8 =>L2Cmd =>L2Sia =>Mpls1Mpls2Mpls3 =>InnerIpv4);
    bins EthMacSec8L2CmdL2SiaMpls1Mpls2Mpls3InnerIpv6Trans = (Eth =>MacSec8 =>L2Cmd =>L2Sia =>Mpls1Mpls2Mpls3 =>InnerIpv6);
    bins EthMacSec8L2CmdL2SiaMpls1Mpls2Mpls3InnerEthTrans = (Eth =>MacSec8 =>L2Cmd =>L2Sia =>Mpls1Mpls2Mpls3 =>InnerEth);
    bins EthMacSec8Tag1qIpv4TcpTrans = (Eth =>MacSec8 =>Tag1q =>Ipv4 =>Tcp);
    bins EthMacSec8Tag1qIpv6TcpTrans = (Eth =>MacSec8 =>Tag1q =>Ipv6 =>Tcp);
    bins EthMacSec8Tag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>Tag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8Tag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>Tag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8Tag1qL2SiaIpv4TcpTrans = (Eth =>MacSec8 =>Tag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec8Tag1qL2SiaIpv6TcpTrans = (Eth =>MacSec8 =>Tag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec8Tag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>Tag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8Tag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>Tag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8Tag1qL2CmdIpv4TcpTrans = (Eth =>MacSec8 =>Tag1q =>L2Cmd =>Ipv4 =>Tcp);
    bins EthMacSec8Tag1qL2CmdIpv6TcpTrans = (Eth =>MacSec8 =>Tag1q =>L2Cmd =>Ipv6 =>Tcp);
    bins EthMacSec8Tag1qL2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8Tag1qL2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8Tag1qL2CmdL2SiaIpv4TcpTrans = (Eth =>MacSec8 =>Tag1q =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec8Tag1qL2CmdL2SiaIpv6TcpTrans = (Eth =>MacSec8 =>Tag1q =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec8Tag1qL2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>Tag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8Tag1qL2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>Tag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8Tag1qTag1qIpv4TcpTrans = (Eth =>MacSec8 =>Tag1qTag1q =>Ipv4 =>Tcp);
    bins EthMacSec8Tag1qTag1qIpv6TcpTrans = (Eth =>MacSec8 =>Tag1qTag1q =>Ipv6 =>Tcp);
    bins EthMacSec8Tag1qTag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>Tag1qTag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8Tag1qTag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>Tag1qTag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8Tag1qTag1qL2SiaIpv4TcpTrans = (Eth =>MacSec8 =>Tag1qTag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec8Tag1qTag1qL2SiaIpv6TcpTrans = (Eth =>MacSec8 =>Tag1qTag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec8Tag1qTag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>Tag1qTag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8Tag1qTag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>Tag1qTag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8Tag1qTag1qL2CmdIpv4TcpTrans = (Eth =>MacSec8 =>Tag1qTag1q =>L2Cmd =>Ipv4 =>Tcp);
    bins EthMacSec8Tag1qTag1qL2CmdIpv6TcpTrans = (Eth =>MacSec8 =>Tag1qTag1q =>L2Cmd =>Ipv6 =>Tcp);
    bins EthMacSec8Tag1qTag1qL2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>Tag1qTag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8Tag1qTag1qL2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>Tag1qTag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8Tag1qTag1qL2CmdL2SiaIpv4TcpTrans = (Eth =>MacSec8 =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec8Tag1qTag1qL2CmdL2SiaIpv6TcpTrans = (Eth =>MacSec8 =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec8Tag1qTag1qL2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8Tag1qTag1qL2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8StagIpv4TcpTrans = (Eth =>MacSec8 =>Stag =>Ipv4 =>Tcp);
    bins EthMacSec8StagIpv6TcpTrans = (Eth =>MacSec8 =>Stag =>Ipv6 =>Tcp);
    bins EthMacSec8StagIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>Stag =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8StagIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>Stag =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8StagL2SiaIpv4TcpTrans = (Eth =>MacSec8 =>Stag =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec8StagL2SiaIpv6TcpTrans = (Eth =>MacSec8 =>Stag =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec8StagL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>Stag =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8StagL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>Stag =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8StagL2CmdIpv4TcpTrans = (Eth =>MacSec8 =>Stag =>L2Cmd =>Ipv4 =>Tcp);
    bins EthMacSec8StagL2CmdIpv6TcpTrans = (Eth =>MacSec8 =>Stag =>L2Cmd =>Ipv6 =>Tcp);
    bins EthMacSec8StagL2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>Stag =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8StagL2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>Stag =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8StagL2CmdL2SiaIpv4TcpTrans = (Eth =>MacSec8 =>Stag =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec8StagL2CmdL2SiaIpv6TcpTrans = (Eth =>MacSec8 =>Stag =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec8StagL2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>Stag =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8StagL2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>Stag =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8StagTag1qIpv4TcpTrans = (Eth =>MacSec8 =>StagTag1q =>Ipv4 =>Tcp);
    bins EthMacSec8StagTag1qIpv6TcpTrans = (Eth =>MacSec8 =>StagTag1q =>Ipv6 =>Tcp);
    bins EthMacSec8StagTag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>StagTag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8StagTag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>StagTag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8StagTag1qL2SiaIpv4TcpTrans = (Eth =>MacSec8 =>StagTag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec8StagTag1qL2SiaIpv6TcpTrans = (Eth =>MacSec8 =>StagTag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec8StagTag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>StagTag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8StagTag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>StagTag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8StagTag1qL2CmdIpv4TcpTrans = (Eth =>MacSec8 =>StagTag1q =>L2Cmd =>Ipv4 =>Tcp);
    bins EthMacSec8StagTag1qL2CmdIpv6TcpTrans = (Eth =>MacSec8 =>StagTag1q =>L2Cmd =>Ipv6 =>Tcp);
    bins EthMacSec8StagTag1qL2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>StagTag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8StagTag1qL2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>StagTag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8StagTag1qL2CmdL2SiaIpv4TcpTrans = (Eth =>MacSec8 =>StagTag1q =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec8StagTag1qL2CmdL2SiaIpv6TcpTrans = (Eth =>MacSec8 =>StagTag1q =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec8StagTag1qL2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>StagTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8StagTag1qL2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>StagTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8VnTagTag1qIpv4TcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1q =>Ipv4 =>Tcp);
    bins EthMacSec8VnTagTag1qIpv6TcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1q =>Ipv6 =>Tcp);
    bins EthMacSec8VnTagTag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8VnTagTag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8VnTagTag1qL2SiaIpv4TcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec8VnTagTag1qL2SiaIpv6TcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec8VnTagTag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8VnTagTag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8VnTagTag1qL2CmdIpv4TcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1q =>L2Cmd =>Ipv4 =>Tcp);
    bins EthMacSec8VnTagTag1qL2CmdIpv6TcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1q =>L2Cmd =>Ipv6 =>Tcp);
    bins EthMacSec8VnTagTag1qL2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8VnTagTag1qL2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8VnTagTag1qL2CmdL2SiaIpv4TcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1q =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec8VnTagTag1qL2CmdL2SiaIpv6TcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1q =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec8VnTagTag1qL2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8VnTagTag1qL2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8VnTagTag1qTag1qIpv4TcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1qTag1q =>Ipv4 =>Tcp);
    bins EthMacSec8VnTagTag1qTag1qIpv6TcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1qTag1q =>Ipv6 =>Tcp);
    bins EthMacSec8VnTagTag1qTag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1qTag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8VnTagTag1qTag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1qTag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8VnTagTag1qTag1qL2SiaIpv4TcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1qTag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec8VnTagTag1qTag1qL2SiaIpv6TcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1qTag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec8VnTagTag1qTag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1qTag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8VnTagTag1qTag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1qTag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8VnTagTag1qTag1qL2CmdIpv4TcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1qTag1q =>L2Cmd =>Ipv4 =>Tcp);
    bins EthMacSec8VnTagTag1qTag1qL2CmdIpv6TcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1qTag1q =>L2Cmd =>Ipv6 =>Tcp);
    bins EthMacSec8VnTagTag1qTag1qL2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1qTag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8VnTagTag1qTag1qL2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1qTag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8VnTagTag1qTag1qL2CmdL2SiaIpv4TcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec8VnTagTag1qTag1qL2CmdL2SiaIpv6TcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec8VnTagTag1qTag1qL2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8VnTagTag1qTag1qL2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>VnTag =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8VnTagStagTag1qIpv4TcpTrans = (Eth =>MacSec8 =>VnTag =>StagTag1q =>Ipv4 =>Tcp);
    bins EthMacSec8VnTagStagTag1qIpv6TcpTrans = (Eth =>MacSec8 =>VnTag =>StagTag1q =>Ipv6 =>Tcp);
    bins EthMacSec8VnTagStagTag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>VnTag =>StagTag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8VnTagStagTag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>VnTag =>StagTag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8VnTagStagTag1qL2SiaIpv4TcpTrans = (Eth =>MacSec8 =>VnTag =>StagTag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec8VnTagStagTag1qL2SiaIpv6TcpTrans = (Eth =>MacSec8 =>VnTag =>StagTag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec8VnTagStagTag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>VnTag =>StagTag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8VnTagStagTag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>VnTag =>StagTag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8VnTagStagTag1qL2CmdIpv4TcpTrans = (Eth =>MacSec8 =>VnTag =>StagTag1q =>L2Cmd =>Ipv4 =>Tcp);
    bins EthMacSec8VnTagStagTag1qL2CmdIpv6TcpTrans = (Eth =>MacSec8 =>VnTag =>StagTag1q =>L2Cmd =>Ipv6 =>Tcp);
    bins EthMacSec8VnTagStagTag1qL2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>VnTag =>StagTag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8VnTagStagTag1qL2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>VnTag =>StagTag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8VnTagStagTag1qL2CmdL2SiaIpv4TcpTrans = (Eth =>MacSec8 =>VnTag =>StagTag1q =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec8VnTagStagTag1qL2CmdL2SiaIpv6TcpTrans = (Eth =>MacSec8 =>VnTag =>StagTag1q =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec8VnTagStagTag1qL2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>VnTag =>StagTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8VnTagStagTag1qL2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>VnTag =>StagTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8SilTag1qIpv4TcpTrans = (Eth =>MacSec8 =>Sil =>Tag1q =>Ipv4 =>Tcp);
    bins EthMacSec8SilTag1qIpv6TcpTrans = (Eth =>MacSec8 =>Sil =>Tag1q =>Ipv6 =>Tcp);
    bins EthMacSec8SilTag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>Sil =>Tag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8SilTag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>Sil =>Tag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8SilTag1qL2SiaIpv4TcpTrans = (Eth =>MacSec8 =>Sil =>Tag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec8SilTag1qL2SiaIpv6TcpTrans = (Eth =>MacSec8 =>Sil =>Tag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec8SilTag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>Sil =>Tag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8SilTag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>Sil =>Tag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8SilTag1qL2CmdIpv4TcpTrans = (Eth =>MacSec8 =>Sil =>Tag1q =>L2Cmd =>Ipv4 =>Tcp);
    bins EthMacSec8SilTag1qL2CmdIpv6TcpTrans = (Eth =>MacSec8 =>Sil =>Tag1q =>L2Cmd =>Ipv6 =>Tcp);
    bins EthMacSec8SilTag1qL2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>Sil =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8SilTag1qL2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>Sil =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8SilTag1qL2CmdL2SiaIpv4TcpTrans = (Eth =>MacSec8 =>Sil =>Tag1q =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec8SilTag1qL2CmdL2SiaIpv6TcpTrans = (Eth =>MacSec8 =>Sil =>Tag1q =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec8SilTag1qL2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>Sil =>Tag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8SilTag1qL2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>Sil =>Tag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8SilTag1qTag1qIpv4TcpTrans = (Eth =>MacSec8 =>Sil =>Tag1qTag1q =>Ipv4 =>Tcp);
    bins EthMacSec8SilTag1qTag1qIpv6TcpTrans = (Eth =>MacSec8 =>Sil =>Tag1qTag1q =>Ipv6 =>Tcp);
    bins EthMacSec8SilTag1qTag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>Sil =>Tag1qTag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8SilTag1qTag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>Sil =>Tag1qTag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8SilTag1qTag1qL2SiaIpv4TcpTrans = (Eth =>MacSec8 =>Sil =>Tag1qTag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec8SilTag1qTag1qL2SiaIpv6TcpTrans = (Eth =>MacSec8 =>Sil =>Tag1qTag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec8SilTag1qTag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>Sil =>Tag1qTag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8SilTag1qTag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>Sil =>Tag1qTag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8SilTag1qTag1qL2CmdIpv4TcpTrans = (Eth =>MacSec8 =>Sil =>Tag1qTag1q =>L2Cmd =>Ipv4 =>Tcp);
    bins EthMacSec8SilTag1qTag1qL2CmdIpv6TcpTrans = (Eth =>MacSec8 =>Sil =>Tag1qTag1q =>L2Cmd =>Ipv6 =>Tcp);
    bins EthMacSec8SilTag1qTag1qL2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>Sil =>Tag1qTag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8SilTag1qTag1qL2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>Sil =>Tag1qTag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8SilTag1qTag1qL2CmdL2SiaIpv4TcpTrans = (Eth =>MacSec8 =>Sil =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec8SilTag1qTag1qL2CmdL2SiaIpv6TcpTrans = (Eth =>MacSec8 =>Sil =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec8SilTag1qTag1qL2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>Sil =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8SilTag1qTag1qL2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>Sil =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8SilVnTagTag1qIpv4TcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1q =>Ipv4 =>Tcp);
    bins EthMacSec8SilVnTagTag1qIpv6TcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1q =>Ipv6 =>Tcp);
    bins EthMacSec8SilVnTagTag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8SilVnTagTag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8SilVnTagTag1qL2SiaIpv4TcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec8SilVnTagTag1qL2SiaIpv6TcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec8SilVnTagTag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8SilVnTagTag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8SilVnTagTag1qL2CmdIpv4TcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1q =>L2Cmd =>Ipv4 =>Tcp);
    bins EthMacSec8SilVnTagTag1qL2CmdIpv6TcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1q =>L2Cmd =>Ipv6 =>Tcp);
    bins EthMacSec8SilVnTagTag1qL2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8SilVnTagTag1qL2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8SilVnTagTag1qL2CmdL2SiaIpv4TcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1q =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec8SilVnTagTag1qL2CmdL2SiaIpv6TcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1q =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec8SilVnTagTag1qL2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8SilVnTagTag1qL2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8SilVnTagTag1qTag1qIpv4TcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1qTag1q =>Ipv4 =>Tcp);
    bins EthMacSec8SilVnTagTag1qTag1qIpv6TcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1qTag1q =>Ipv6 =>Tcp);
    bins EthMacSec8SilVnTagTag1qTag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1qTag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8SilVnTagTag1qTag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1qTag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8SilVnTagTag1qTag1qL2SiaIpv4TcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1qTag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec8SilVnTagTag1qTag1qL2SiaIpv6TcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1qTag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec8SilVnTagTag1qTag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1qTag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8SilVnTagTag1qTag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1qTag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8SilVnTagTag1qTag1qL2CmdIpv4TcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1qTag1q =>L2Cmd =>Ipv4 =>Tcp);
    bins EthMacSec8SilVnTagTag1qTag1qL2CmdIpv6TcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1qTag1q =>L2Cmd =>Ipv6 =>Tcp);
    bins EthMacSec8SilVnTagTag1qTag1qL2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1qTag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8SilVnTagTag1qTag1qL2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1qTag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec8SilVnTagTag1qTag1qL2CmdL2SiaIpv4TcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec8SilVnTagTag1qTag1qL2CmdL2SiaIpv6TcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec8SilVnTagTag1qTag1qL2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec8SilVnTagTag1qTag1qL2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec8 =>Sil =>VnTag =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16Ipv4TcpTrans = (Eth =>MacSec16 =>Ipv4 =>Tcp);
    bins EthMacSec16Ipv6TcpTrans = (Eth =>MacSec16 =>Ipv6 =>Tcp);
    bins EthMacSec16Ipv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16Ipv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16Mpls1InnerIpv4Trans = (Eth =>MacSec16 =>Mpls1 =>InnerIpv4);
    bins EthMacSec16Mpls1InnerIpv6Trans = (Eth =>MacSec16 =>Mpls1 =>InnerIpv6);
    bins EthMacSec16Mpls1InnerEthTrans = (Eth =>MacSec16 =>Mpls1 =>InnerEth);
    bins EthMacSec16Mpls1Mpls2InnerIpv4Trans = (Eth =>MacSec16 =>Mpls1Mpls2 =>InnerIpv4);
    bins EthMacSec16Mpls1Mpls2InnerIpv6Trans = (Eth =>MacSec16 =>Mpls1Mpls2 =>InnerIpv6);
    bins EthMacSec16Mpls1Mpls2InnerEthTrans = (Eth =>MacSec16 =>Mpls1Mpls2 =>InnerEth);
    bins EthMacSec16Mpls1Mpls2Mpls3InnerIpv4Trans = (Eth =>MacSec16 =>Mpls1Mpls2Mpls3 =>InnerIpv4);
    bins EthMacSec16Mpls1Mpls2Mpls3InnerIpv6Trans = (Eth =>MacSec16 =>Mpls1Mpls2Mpls3 =>InnerIpv6);
    bins EthMacSec16Mpls1Mpls2Mpls3InnerEthTrans = (Eth =>MacSec16 =>Mpls1Mpls2Mpls3 =>InnerEth);
    bins EthMacSec16L2SiaIpv4TcpTrans = (Eth =>MacSec16 =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec16L2SiaIpv6TcpTrans = (Eth =>MacSec16 =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec16L2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16L2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16L2SiaMpls1InnerIpv4Trans = (Eth =>MacSec16 =>L2Sia =>Mpls1 =>InnerIpv4);
    bins EthMacSec16L2SiaMpls1InnerIpv6Trans = (Eth =>MacSec16 =>L2Sia =>Mpls1 =>InnerIpv6);
    bins EthMacSec16L2SiaMpls1InnerEthTrans = (Eth =>MacSec16 =>L2Sia =>Mpls1 =>InnerEth);
    bins EthMacSec16L2SiaMpls1Mpls2InnerIpv4Trans = (Eth =>MacSec16 =>L2Sia =>Mpls1Mpls2 =>InnerIpv4);
    bins EthMacSec16L2SiaMpls1Mpls2InnerIpv6Trans = (Eth =>MacSec16 =>L2Sia =>Mpls1Mpls2 =>InnerIpv6);
    bins EthMacSec16L2SiaMpls1Mpls2InnerEthTrans = (Eth =>MacSec16 =>L2Sia =>Mpls1Mpls2 =>InnerEth);
    bins EthMacSec16L2SiaMpls1Mpls2Mpls3InnerIpv4Trans = (Eth =>MacSec16 =>L2Sia =>Mpls1Mpls2Mpls3 =>InnerIpv4);
    bins EthMacSec16L2SiaMpls1Mpls2Mpls3InnerIpv6Trans = (Eth =>MacSec16 =>L2Sia =>Mpls1Mpls2Mpls3 =>InnerIpv6);
    bins EthMacSec16L2SiaMpls1Mpls2Mpls3InnerEthTrans = (Eth =>MacSec16 =>L2Sia =>Mpls1Mpls2Mpls3 =>InnerEth);
    bins EthMacSec16L2CmdIpv4TcpTrans = (Eth =>MacSec16 =>L2Cmd =>Ipv4 =>Tcp);
    bins EthMacSec16L2CmdIpv6TcpTrans = (Eth =>MacSec16 =>L2Cmd =>Ipv6 =>Tcp);
    bins EthMacSec16L2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16L2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16L2CmdMpls1InnerIpv4Trans = (Eth =>MacSec16 =>L2Cmd =>Mpls1 =>InnerIpv4);
    bins EthMacSec16L2CmdMpls1InnerIpv6Trans = (Eth =>MacSec16 =>L2Cmd =>Mpls1 =>InnerIpv6);
    bins EthMacSec16L2CmdMpls1InnerEthTrans = (Eth =>MacSec16 =>L2Cmd =>Mpls1 =>InnerEth);
    bins EthMacSec16L2CmdMpls1Mpls2InnerIpv4Trans = (Eth =>MacSec16 =>L2Cmd =>Mpls1Mpls2 =>InnerIpv4);
    bins EthMacSec16L2CmdMpls1Mpls2InnerIpv6Trans = (Eth =>MacSec16 =>L2Cmd =>Mpls1Mpls2 =>InnerIpv6);
    bins EthMacSec16L2CmdMpls1Mpls2InnerEthTrans = (Eth =>MacSec16 =>L2Cmd =>Mpls1Mpls2 =>InnerEth);
    bins EthMacSec16L2CmdMpls1Mpls2Mpls3InnerIpv4Trans = (Eth =>MacSec16 =>L2Cmd =>Mpls1Mpls2Mpls3 =>InnerIpv4);
    bins EthMacSec16L2CmdMpls1Mpls2Mpls3InnerIpv6Trans = (Eth =>MacSec16 =>L2Cmd =>Mpls1Mpls2Mpls3 =>InnerIpv6);
    bins EthMacSec16L2CmdMpls1Mpls2Mpls3InnerEthTrans = (Eth =>MacSec16 =>L2Cmd =>Mpls1Mpls2Mpls3 =>InnerEth);
    bins EthMacSec16L2CmdL2SiaIpv4TcpTrans = (Eth =>MacSec16 =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec16L2CmdL2SiaIpv6TcpTrans = (Eth =>MacSec16 =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec16L2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16L2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16L2CmdL2SiaMpls1InnerIpv4Trans = (Eth =>MacSec16 =>L2Cmd =>L2Sia =>Mpls1 =>InnerIpv4);
    bins EthMacSec16L2CmdL2SiaMpls1InnerIpv6Trans = (Eth =>MacSec16 =>L2Cmd =>L2Sia =>Mpls1 =>InnerIpv6);
    bins EthMacSec16L2CmdL2SiaMpls1InnerEthTrans = (Eth =>MacSec16 =>L2Cmd =>L2Sia =>Mpls1 =>InnerEth);
    bins EthMacSec16L2CmdL2SiaMpls1Mpls2InnerIpv4Trans = (Eth =>MacSec16 =>L2Cmd =>L2Sia =>Mpls1Mpls2 =>InnerIpv4);
    bins EthMacSec16L2CmdL2SiaMpls1Mpls2InnerIpv6Trans = (Eth =>MacSec16 =>L2Cmd =>L2Sia =>Mpls1Mpls2 =>InnerIpv6);
    bins EthMacSec16L2CmdL2SiaMpls1Mpls2InnerEthTrans = (Eth =>MacSec16 =>L2Cmd =>L2Sia =>Mpls1Mpls2 =>InnerEth);
    bins EthMacSec16L2CmdL2SiaMpls1Mpls2Mpls3InnerIpv4Trans = (Eth =>MacSec16 =>L2Cmd =>L2Sia =>Mpls1Mpls2Mpls3 =>InnerIpv4);
    bins EthMacSec16L2CmdL2SiaMpls1Mpls2Mpls3InnerIpv6Trans = (Eth =>MacSec16 =>L2Cmd =>L2Sia =>Mpls1Mpls2Mpls3 =>InnerIpv6);
    bins EthMacSec16L2CmdL2SiaMpls1Mpls2Mpls3InnerEthTrans = (Eth =>MacSec16 =>L2Cmd =>L2Sia =>Mpls1Mpls2Mpls3 =>InnerEth);
    bins EthMacSec16Tag1qIpv4TcpTrans = (Eth =>MacSec16 =>Tag1q =>Ipv4 =>Tcp);
    bins EthMacSec16Tag1qIpv6TcpTrans = (Eth =>MacSec16 =>Tag1q =>Ipv6 =>Tcp);
    bins EthMacSec16Tag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>Tag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16Tag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>Tag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16Tag1qL2SiaIpv4TcpTrans = (Eth =>MacSec16 =>Tag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec16Tag1qL2SiaIpv6TcpTrans = (Eth =>MacSec16 =>Tag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec16Tag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>Tag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16Tag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>Tag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16Tag1qL2CmdIpv4TcpTrans = (Eth =>MacSec16 =>Tag1q =>L2Cmd =>Ipv4 =>Tcp);
    bins EthMacSec16Tag1qL2CmdIpv6TcpTrans = (Eth =>MacSec16 =>Tag1q =>L2Cmd =>Ipv6 =>Tcp);
    bins EthMacSec16Tag1qL2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16Tag1qL2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16Tag1qL2CmdL2SiaIpv4TcpTrans = (Eth =>MacSec16 =>Tag1q =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec16Tag1qL2CmdL2SiaIpv6TcpTrans = (Eth =>MacSec16 =>Tag1q =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec16Tag1qL2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>Tag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16Tag1qL2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>Tag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16Tag1qTag1qIpv4TcpTrans = (Eth =>MacSec16 =>Tag1qTag1q =>Ipv4 =>Tcp);
    bins EthMacSec16Tag1qTag1qIpv6TcpTrans = (Eth =>MacSec16 =>Tag1qTag1q =>Ipv6 =>Tcp);
    bins EthMacSec16Tag1qTag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>Tag1qTag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16Tag1qTag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>Tag1qTag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16Tag1qTag1qL2SiaIpv4TcpTrans = (Eth =>MacSec16 =>Tag1qTag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec16Tag1qTag1qL2SiaIpv6TcpTrans = (Eth =>MacSec16 =>Tag1qTag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec16Tag1qTag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>Tag1qTag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16Tag1qTag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>Tag1qTag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16Tag1qTag1qL2CmdIpv4TcpTrans = (Eth =>MacSec16 =>Tag1qTag1q =>L2Cmd =>Ipv4 =>Tcp);
    bins EthMacSec16Tag1qTag1qL2CmdIpv6TcpTrans = (Eth =>MacSec16 =>Tag1qTag1q =>L2Cmd =>Ipv6 =>Tcp);
    bins EthMacSec16Tag1qTag1qL2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>Tag1qTag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16Tag1qTag1qL2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>Tag1qTag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16Tag1qTag1qL2CmdL2SiaIpv4TcpTrans = (Eth =>MacSec16 =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec16Tag1qTag1qL2CmdL2SiaIpv6TcpTrans = (Eth =>MacSec16 =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec16Tag1qTag1qL2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16Tag1qTag1qL2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16StagIpv4TcpTrans = (Eth =>MacSec16 =>Stag =>Ipv4 =>Tcp);
    bins EthMacSec16StagIpv6TcpTrans = (Eth =>MacSec16 =>Stag =>Ipv6 =>Tcp);
    bins EthMacSec16StagIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>Stag =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16StagIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>Stag =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16StagL2SiaIpv4TcpTrans = (Eth =>MacSec16 =>Stag =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec16StagL2SiaIpv6TcpTrans = (Eth =>MacSec16 =>Stag =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec16StagL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>Stag =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16StagL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>Stag =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16StagL2CmdIpv4TcpTrans = (Eth =>MacSec16 =>Stag =>L2Cmd =>Ipv4 =>Tcp);
    bins EthMacSec16StagL2CmdIpv6TcpTrans = (Eth =>MacSec16 =>Stag =>L2Cmd =>Ipv6 =>Tcp);
    bins EthMacSec16StagL2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>Stag =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16StagL2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>Stag =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16StagL2CmdL2SiaIpv4TcpTrans = (Eth =>MacSec16 =>Stag =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec16StagL2CmdL2SiaIpv6TcpTrans = (Eth =>MacSec16 =>Stag =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec16StagL2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>Stag =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16StagL2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>Stag =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16StagTag1qIpv4TcpTrans = (Eth =>MacSec16 =>StagTag1q =>Ipv4 =>Tcp);
    bins EthMacSec16StagTag1qIpv6TcpTrans = (Eth =>MacSec16 =>StagTag1q =>Ipv6 =>Tcp);
    bins EthMacSec16StagTag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>StagTag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16StagTag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>StagTag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16StagTag1qL2SiaIpv4TcpTrans = (Eth =>MacSec16 =>StagTag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec16StagTag1qL2SiaIpv6TcpTrans = (Eth =>MacSec16 =>StagTag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec16StagTag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>StagTag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16StagTag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>StagTag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16StagTag1qL2CmdIpv4TcpTrans = (Eth =>MacSec16 =>StagTag1q =>L2Cmd =>Ipv4 =>Tcp);
    bins EthMacSec16StagTag1qL2CmdIpv6TcpTrans = (Eth =>MacSec16 =>StagTag1q =>L2Cmd =>Ipv6 =>Tcp);
    bins EthMacSec16StagTag1qL2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>StagTag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16StagTag1qL2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>StagTag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16StagTag1qL2CmdL2SiaIpv4TcpTrans = (Eth =>MacSec16 =>StagTag1q =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec16StagTag1qL2CmdL2SiaIpv6TcpTrans = (Eth =>MacSec16 =>StagTag1q =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec16StagTag1qL2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>StagTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16StagTag1qL2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>StagTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16VnTagTag1qIpv4TcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1q =>Ipv4 =>Tcp);
    bins EthMacSec16VnTagTag1qIpv6TcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1q =>Ipv6 =>Tcp);
    bins EthMacSec16VnTagTag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16VnTagTag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16VnTagTag1qL2SiaIpv4TcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec16VnTagTag1qL2SiaIpv6TcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec16VnTagTag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16VnTagTag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16VnTagTag1qL2CmdIpv4TcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1q =>L2Cmd =>Ipv4 =>Tcp);
    bins EthMacSec16VnTagTag1qL2CmdIpv6TcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1q =>L2Cmd =>Ipv6 =>Tcp);
    bins EthMacSec16VnTagTag1qL2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16VnTagTag1qL2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16VnTagTag1qL2CmdL2SiaIpv4TcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1q =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec16VnTagTag1qL2CmdL2SiaIpv6TcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1q =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec16VnTagTag1qL2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16VnTagTag1qL2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16VnTagTag1qTag1qIpv4TcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1qTag1q =>Ipv4 =>Tcp);
    bins EthMacSec16VnTagTag1qTag1qIpv6TcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1qTag1q =>Ipv6 =>Tcp);
    bins EthMacSec16VnTagTag1qTag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1qTag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16VnTagTag1qTag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1qTag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16VnTagTag1qTag1qL2SiaIpv4TcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1qTag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec16VnTagTag1qTag1qL2SiaIpv6TcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1qTag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec16VnTagTag1qTag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1qTag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16VnTagTag1qTag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1qTag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16VnTagTag1qTag1qL2CmdIpv4TcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1qTag1q =>L2Cmd =>Ipv4 =>Tcp);
    bins EthMacSec16VnTagTag1qTag1qL2CmdIpv6TcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1qTag1q =>L2Cmd =>Ipv6 =>Tcp);
    bins EthMacSec16VnTagTag1qTag1qL2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1qTag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16VnTagTag1qTag1qL2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1qTag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16VnTagTag1qTag1qL2CmdL2SiaIpv4TcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec16VnTagTag1qTag1qL2CmdL2SiaIpv6TcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec16VnTagTag1qTag1qL2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16VnTagTag1qTag1qL2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>VnTag =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16VnTagStagTag1qIpv4TcpTrans = (Eth =>MacSec16 =>VnTag =>StagTag1q =>Ipv4 =>Tcp);
    bins EthMacSec16VnTagStagTag1qIpv6TcpTrans = (Eth =>MacSec16 =>VnTag =>StagTag1q =>Ipv6 =>Tcp);
    bins EthMacSec16VnTagStagTag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>VnTag =>StagTag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16VnTagStagTag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>VnTag =>StagTag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16VnTagStagTag1qL2SiaIpv4TcpTrans = (Eth =>MacSec16 =>VnTag =>StagTag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec16VnTagStagTag1qL2SiaIpv6TcpTrans = (Eth =>MacSec16 =>VnTag =>StagTag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec16VnTagStagTag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>VnTag =>StagTag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16VnTagStagTag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>VnTag =>StagTag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16VnTagStagTag1qL2CmdIpv4TcpTrans = (Eth =>MacSec16 =>VnTag =>StagTag1q =>L2Cmd =>Ipv4 =>Tcp);
    bins EthMacSec16VnTagStagTag1qL2CmdIpv6TcpTrans = (Eth =>MacSec16 =>VnTag =>StagTag1q =>L2Cmd =>Ipv6 =>Tcp);
    bins EthMacSec16VnTagStagTag1qL2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>VnTag =>StagTag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16VnTagStagTag1qL2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>VnTag =>StagTag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16VnTagStagTag1qL2CmdL2SiaIpv4TcpTrans = (Eth =>MacSec16 =>VnTag =>StagTag1q =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec16VnTagStagTag1qL2CmdL2SiaIpv6TcpTrans = (Eth =>MacSec16 =>VnTag =>StagTag1q =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec16VnTagStagTag1qL2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>VnTag =>StagTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16VnTagStagTag1qL2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>VnTag =>StagTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16SilTag1qIpv4TcpTrans = (Eth =>MacSec16 =>Sil =>Tag1q =>Ipv4 =>Tcp);
    bins EthMacSec16SilTag1qIpv6TcpTrans = (Eth =>MacSec16 =>Sil =>Tag1q =>Ipv6 =>Tcp);
    bins EthMacSec16SilTag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>Sil =>Tag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16SilTag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>Sil =>Tag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16SilTag1qL2SiaIpv4TcpTrans = (Eth =>MacSec16 =>Sil =>Tag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec16SilTag1qL2SiaIpv6TcpTrans = (Eth =>MacSec16 =>Sil =>Tag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec16SilTag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>Sil =>Tag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16SilTag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>Sil =>Tag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16SilTag1qL2CmdIpv4TcpTrans = (Eth =>MacSec16 =>Sil =>Tag1q =>L2Cmd =>Ipv4 =>Tcp);
    bins EthMacSec16SilTag1qL2CmdIpv6TcpTrans = (Eth =>MacSec16 =>Sil =>Tag1q =>L2Cmd =>Ipv6 =>Tcp);
    bins EthMacSec16SilTag1qL2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>Sil =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16SilTag1qL2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>Sil =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16SilTag1qL2CmdL2SiaIpv4TcpTrans = (Eth =>MacSec16 =>Sil =>Tag1q =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec16SilTag1qL2CmdL2SiaIpv6TcpTrans = (Eth =>MacSec16 =>Sil =>Tag1q =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec16SilTag1qL2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>Sil =>Tag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16SilTag1qL2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>Sil =>Tag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16SilTag1qTag1qIpv4TcpTrans = (Eth =>MacSec16 =>Sil =>Tag1qTag1q =>Ipv4 =>Tcp);
    bins EthMacSec16SilTag1qTag1qIpv6TcpTrans = (Eth =>MacSec16 =>Sil =>Tag1qTag1q =>Ipv6 =>Tcp);
    bins EthMacSec16SilTag1qTag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>Sil =>Tag1qTag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16SilTag1qTag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>Sil =>Tag1qTag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16SilTag1qTag1qL2SiaIpv4TcpTrans = (Eth =>MacSec16 =>Sil =>Tag1qTag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec16SilTag1qTag1qL2SiaIpv6TcpTrans = (Eth =>MacSec16 =>Sil =>Tag1qTag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec16SilTag1qTag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>Sil =>Tag1qTag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16SilTag1qTag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>Sil =>Tag1qTag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16SilTag1qTag1qL2CmdIpv4TcpTrans = (Eth =>MacSec16 =>Sil =>Tag1qTag1q =>L2Cmd =>Ipv4 =>Tcp);
    bins EthMacSec16SilTag1qTag1qL2CmdIpv6TcpTrans = (Eth =>MacSec16 =>Sil =>Tag1qTag1q =>L2Cmd =>Ipv6 =>Tcp);
    bins EthMacSec16SilTag1qTag1qL2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>Sil =>Tag1qTag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16SilTag1qTag1qL2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>Sil =>Tag1qTag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16SilTag1qTag1qL2CmdL2SiaIpv4TcpTrans = (Eth =>MacSec16 =>Sil =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec16SilTag1qTag1qL2CmdL2SiaIpv6TcpTrans = (Eth =>MacSec16 =>Sil =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec16SilTag1qTag1qL2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>Sil =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16SilTag1qTag1qL2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>Sil =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16SilVnTagTag1qIpv4TcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1q =>Ipv4 =>Tcp);
    bins EthMacSec16SilVnTagTag1qIpv6TcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1q =>Ipv6 =>Tcp);
    bins EthMacSec16SilVnTagTag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16SilVnTagTag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16SilVnTagTag1qL2SiaIpv4TcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec16SilVnTagTag1qL2SiaIpv6TcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec16SilVnTagTag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16SilVnTagTag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16SilVnTagTag1qL2CmdIpv4TcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1q =>L2Cmd =>Ipv4 =>Tcp);
    bins EthMacSec16SilVnTagTag1qL2CmdIpv6TcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1q =>L2Cmd =>Ipv6 =>Tcp);
    bins EthMacSec16SilVnTagTag1qL2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16SilVnTagTag1qL2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16SilVnTagTag1qL2CmdL2SiaIpv4TcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1q =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec16SilVnTagTag1qL2CmdL2SiaIpv6TcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1q =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec16SilVnTagTag1qL2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16SilVnTagTag1qL2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16SilVnTagTag1qTag1qIpv4TcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1qTag1q =>Ipv4 =>Tcp);
    bins EthMacSec16SilVnTagTag1qTag1qIpv6TcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1qTag1q =>Ipv6 =>Tcp);
    bins EthMacSec16SilVnTagTag1qTag1qIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1qTag1q =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16SilVnTagTag1qTag1qIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1qTag1q =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16SilVnTagTag1qTag1qL2SiaIpv4TcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1qTag1q =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec16SilVnTagTag1qTag1qL2SiaIpv6TcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1qTag1q =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec16SilVnTagTag1qTag1qL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1qTag1q =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16SilVnTagTag1qTag1qL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1qTag1q =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16SilVnTagTag1qTag1qL2CmdIpv4TcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1qTag1q =>L2Cmd =>Ipv4 =>Tcp);
    bins EthMacSec16SilVnTagTag1qTag1qL2CmdIpv6TcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1qTag1q =>L2Cmd =>Ipv6 =>Tcp);
    bins EthMacSec16SilVnTagTag1qTag1qL2CmdIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1qTag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16SilVnTagTag1qTag1qL2CmdIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1qTag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthMacSec16SilVnTagTag1qTag1qL2CmdL2SiaIpv4TcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv4 =>Tcp);
    bins EthMacSec16SilVnTagTag1qTag1qL2CmdL2SiaIpv6TcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6 =>Tcp);
    bins EthMacSec16SilVnTagTag1qTag1qL2CmdL2SiaIpv6Ipv6ExtnDstnOption2TcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnDstnOption2 =>Tcp);
    bins EthMacSec16SilVnTagTag1qTag1qL2CmdL2SiaIpv6Ipv6ExtnFragmentTcpTrans = (Eth =>MacSec16 =>Sil =>VnTag =>Tag1qTag1q =>L2Cmd =>L2Sia =>Ipv6Ipv6ExtnFragment =>Tcp);
    bins EthArpTrans = (Eth =>Arp);
    bins EthRarpTrans = (Eth =>Rarp);
    bins EthTag1qArpTrans = (Eth =>Tag1q =>Arp);
    bins EthTag1qRarpTrans = (Eth =>Tag1q =>Rarp);
    bins EthVnTagTag1qArpTrans = (Eth =>VnTag =>Tag1q =>Arp);
    bins EthVnTagTag1qRarpTrans = (Eth =>VnTag =>Tag1q =>Rarp);
    bins EthVnTagTag1qL2CmdArpTrans = (Eth =>VnTag =>Tag1q =>L2Cmd =>Arp);
    bins EthVnTagTag1qL2CmdRarpTrans = (Eth =>VnTag =>Tag1q =>L2Cmd =>Rarp);
    bins EthMacSec8ArpTrans = (Eth =>MacSec8 =>Arp);
    bins EthMacSec8RarpTrans = (Eth =>MacSec8 =>Rarp);
    bins EthMacSec8L2CmdArpTrans = (Eth =>MacSec8 =>L2Cmd =>Arp);
    bins EthMacSec8L2CmdRarpTrans = (Eth =>MacSec8 =>L2Cmd =>Rarp);
    bins EthMacSec8Tag1qArpTrans = (Eth =>MacSec8 =>Tag1q =>Arp);
    bins EthMacSec8Tag1qRarpTrans = (Eth =>MacSec8 =>Tag1q =>Rarp);
    bins EthMacSec8Tag1qL2CmdArpTrans = (Eth =>MacSec8 =>Tag1q =>L2Cmd =>Arp);
    bins EthMacSec8Tag1qL2CmdRarpTrans = (Eth =>MacSec8 =>Tag1q =>L2Cmd =>Rarp);
    bins EthMacSec8VnTagTag1qArpTrans = (Eth =>MacSec8 =>VnTag =>Tag1q =>Arp);
    bins EthMacSec8VnTagTag1qRarpTrans = (Eth =>MacSec8 =>VnTag =>Tag1q =>Rarp);
    bins EthMacSec8VnTagTag1qL2CmdArpTrans = (Eth =>MacSec8 =>VnTag =>Tag1q =>L2Cmd =>Arp);
    bins EthMacSec8VnTagTag1qL2CmdRarpTrans = (Eth =>MacSec8 =>VnTag =>Tag1q =>L2Cmd =>Rarp);
    bins EthMacSec16ArpTrans = (Eth =>MacSec16 =>Arp);
    bins EthMacSec16RarpTrans = (Eth =>MacSec16 =>Rarp);
    bins EthMacSec16L2CmdArpTrans = (Eth =>MacSec16 =>L2Cmd =>Arp);
    bins EthMacSec16L2CmdRarpTrans = (Eth =>MacSec16 =>L2Cmd =>Rarp);
    bins EthMacSec16Tag1qArpTrans = (Eth =>MacSec16 =>Tag1q =>Arp);
    bins EthMacSec16Tag1qRarpTrans = (Eth =>MacSec16 =>Tag1q =>Rarp);
    bins EthMacSec16Tag1qL2CmdArpTrans = (Eth =>MacSec16 =>Tag1q =>L2Cmd =>Arp);
    bins EthMacSec16Tag1qL2CmdRarpTrans = (Eth =>MacSec16 =>Tag1q =>L2Cmd =>Rarp);
    bins EthMacSec16VnTagTag1qArpTrans = (Eth =>MacSec16 =>VnTag =>Tag1q =>Arp);
    bins EthMacSec16VnTagTag1qRarpTrans = (Eth =>MacSec16 =>VnTag =>Tag1q =>Rarp);
    bins EthMacSec16VnTagTag1qL2CmdArpTrans = (Eth =>MacSec16 =>VnTag =>Tag1q =>L2Cmd =>Arp);
    bins EthMacSec16VnTagTag1qL2CmdRarpTrans = (Eth =>MacSec16 =>VnTag =>Tag1q =>L2Cmd =>Rarp);
    bins EthL2_1588Trans = (Eth =>L2_1588);
    bins EthTag1qL2_1588Trans = (Eth =>Tag1q =>L2_1588);
    bins EthVnTagTag1qL2_1588Trans = (Eth =>VnTag =>Tag1q =>L2_1588);
    bins EthVnTagTag1qL2CmdL2_1588Trans = (Eth =>VnTag =>Tag1q =>L2Cmd =>L2_1588);
    bins EthMacSec8L2_1588Trans = (Eth =>MacSec8 =>L2_1588);
    bins EthMacSec8L2CmdL2_1588Trans = (Eth =>MacSec8 =>L2Cmd =>L2_1588);
    bins EthMacSec8Tag1qL2_1588Trans = (Eth =>MacSec8 =>Tag1q =>L2_1588);
    bins EthMacSec8Tag1qL2CmdL2_1588Trans = (Eth =>MacSec8 =>Tag1q =>L2Cmd =>L2_1588);
    bins EthMacSec8VnTagTag1qL2_1588Trans = (Eth =>MacSec8 =>VnTag =>Tag1q =>L2_1588);
    bins EthMacSec8VnTagTag1qL2CmdL2_1588Trans = (Eth =>MacSec8 =>VnTag =>Tag1q =>L2Cmd =>L2_1588);
    bins EthMacSec16L2_1588Trans = (Eth =>MacSec16 =>L2_1588);
    bins EthMacSec16L2CmdL2_1588Trans = (Eth =>MacSec16 =>L2Cmd =>L2_1588);
    bins EthMacSec16Tag1qL2_1588Trans = (Eth =>MacSec16 =>Tag1q =>L2_1588);
    bins EthMacSec16Tag1qL2CmdL2_1588Trans = (Eth =>MacSec16 =>Tag1q =>L2Cmd =>L2_1588);
    bins EthMacSec16VnTagTag1qL2_1588Trans = (Eth =>MacSec16 =>VnTag =>Tag1q =>L2_1588);
    bins EthMacSec16VnTagTag1qL2CmdL2_1588Trans = (Eth =>MacSec16 =>VnTag =>Tag1q =>L2Cmd =>L2_1588);
    bins EthIpv4UdpL3_1588Trans = (Eth =>Ipv4 =>Udp =>L3_1588);
    bins EthIpv6UdpL3_1588Trans = (Eth =>Ipv6 =>Udp =>L3_1588);
    bins EthIpv6Ipv6ExtnDstnOption2UdpL3_1588Trans = (Eth =>Ipv6Ipv6ExtnDstnOption2 =>Udp =>L3_1588);
    bins EthIpv6Ipv6ExtnFragmentUdpL3_1588Trans = (Eth =>Ipv6Ipv6ExtnFragment =>Udp =>L3_1588);
    bins EthTag1qIpv4UdpL3_1588Trans = (Eth =>Tag1q =>Ipv4 =>Udp =>L3_1588);
    bins EthTag1qIpv6UdpL3_1588Trans = (Eth =>Tag1q =>Ipv6 =>Udp =>L3_1588);
    bins EthTag1qIpv6Ipv6ExtnDstnOption2UdpL3_1588Trans = (Eth =>Tag1q =>Ipv6Ipv6ExtnDstnOption2 =>Udp =>L3_1588);
    bins EthTag1qIpv6Ipv6ExtnFragmentUdpL3_1588Trans = (Eth =>Tag1q =>Ipv6Ipv6ExtnFragment =>Udp =>L3_1588);
    bins EthVnTagTag1qIpv4UdpL3_1588Trans = (Eth =>VnTag =>Tag1q =>Ipv4 =>Udp =>L3_1588);
    bins EthVnTagTag1qIpv6UdpL3_1588Trans = (Eth =>VnTag =>Tag1q =>Ipv6 =>Udp =>L3_1588);
    bins EthVnTagTag1qIpv6Ipv6ExtnDstnOption2UdpL3_1588Trans = (Eth =>VnTag =>Tag1q =>Ipv6Ipv6ExtnDstnOption2 =>Udp =>L3_1588);
    bins EthVnTagTag1qIpv6Ipv6ExtnFragmentUdpL3_1588Trans = (Eth =>VnTag =>Tag1q =>Ipv6Ipv6ExtnFragment =>Udp =>L3_1588);
    bins EthVnTagTag1qL2CmdIpv4UdpL3_1588Trans = (Eth =>VnTag =>Tag1q =>L2Cmd =>Ipv4 =>Udp =>L3_1588);
    bins EthVnTagTag1qL2CmdIpv6UdpL3_1588Trans = (Eth =>VnTag =>Tag1q =>L2Cmd =>Ipv6 =>Udp =>L3_1588);
    bins EthVnTagTag1qL2CmdIpv6Ipv6ExtnDstnOption2UdpL3_1588Trans = (Eth =>VnTag =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Udp =>L3_1588);
    bins EthVnTagTag1qL2CmdIpv6Ipv6ExtnFragmentUdpL3_1588Trans = (Eth =>VnTag =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Udp =>L3_1588);
    bins EthMacSec8Ipv4UdpL3_1588Trans = (Eth =>MacSec8 =>Ipv4 =>Udp =>L3_1588);
    bins EthMacSec8Ipv6UdpL3_1588Trans = (Eth =>MacSec8 =>Ipv6 =>Udp =>L3_1588);
    bins EthMacSec8Ipv6Ipv6ExtnDstnOption2UdpL3_1588Trans = (Eth =>MacSec8 =>Ipv6Ipv6ExtnDstnOption2 =>Udp =>L3_1588);
    bins EthMacSec8Ipv6Ipv6ExtnFragmentUdpL3_1588Trans = (Eth =>MacSec8 =>Ipv6Ipv6ExtnFragment =>Udp =>L3_1588);
    bins EthMacSec8L2CmdIpv4UdpL3_1588Trans = (Eth =>MacSec8 =>L2Cmd =>Ipv4 =>Udp =>L3_1588);
    bins EthMacSec8L2CmdIpv6UdpL3_1588Trans = (Eth =>MacSec8 =>L2Cmd =>Ipv6 =>Udp =>L3_1588);
    bins EthMacSec8L2CmdIpv6Ipv6ExtnDstnOption2UdpL3_1588Trans = (Eth =>MacSec8 =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Udp =>L3_1588);
    bins EthMacSec8L2CmdIpv6Ipv6ExtnFragmentUdpL3_1588Trans = (Eth =>MacSec8 =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Udp =>L3_1588);
    bins EthMacSec8Tag1qIpv4UdpL3_1588Trans = (Eth =>MacSec8 =>Tag1q =>Ipv4 =>Udp =>L3_1588);
    bins EthMacSec8Tag1qIpv6UdpL3_1588Trans = (Eth =>MacSec8 =>Tag1q =>Ipv6 =>Udp =>L3_1588);
    bins EthMacSec8Tag1qIpv6Ipv6ExtnDstnOption2UdpL3_1588Trans = (Eth =>MacSec8 =>Tag1q =>Ipv6Ipv6ExtnDstnOption2 =>Udp =>L3_1588);
    bins EthMacSec8Tag1qIpv6Ipv6ExtnFragmentUdpL3_1588Trans = (Eth =>MacSec8 =>Tag1q =>Ipv6Ipv6ExtnFragment =>Udp =>L3_1588);
    bins EthMacSec8Tag1qL2CmdIpv4UdpL3_1588Trans = (Eth =>MacSec8 =>Tag1q =>L2Cmd =>Ipv4 =>Udp =>L3_1588);
    bins EthMacSec8Tag1qL2CmdIpv6UdpL3_1588Trans = (Eth =>MacSec8 =>Tag1q =>L2Cmd =>Ipv6 =>Udp =>L3_1588);
    bins EthMacSec8Tag1qL2CmdIpv6Ipv6ExtnDstnOption2UdpL3_1588Trans = (Eth =>MacSec8 =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Udp =>L3_1588);
    bins EthMacSec8Tag1qL2CmdIpv6Ipv6ExtnFragmentUdpL3_1588Trans = (Eth =>MacSec8 =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Udp =>L3_1588);
    bins EthMacSec8VnTagTag1qIpv4UdpL3_1588Trans = (Eth =>MacSec8 =>VnTag =>Tag1q =>Ipv4 =>Udp =>L3_1588);
    bins EthMacSec8VnTagTag1qIpv6UdpL3_1588Trans = (Eth =>MacSec8 =>VnTag =>Tag1q =>Ipv6 =>Udp =>L3_1588);
    bins EthMacSec8VnTagTag1qIpv6Ipv6ExtnDstnOption2UdpL3_1588Trans = (Eth =>MacSec8 =>VnTag =>Tag1q =>Ipv6Ipv6ExtnDstnOption2 =>Udp =>L3_1588);
    bins EthMacSec8VnTagTag1qIpv6Ipv6ExtnFragmentUdpL3_1588Trans = (Eth =>MacSec8 =>VnTag =>Tag1q =>Ipv6Ipv6ExtnFragment =>Udp =>L3_1588);
    bins EthMacSec8VnTagTag1qL2CmdIpv4UdpL3_1588Trans = (Eth =>MacSec8 =>VnTag =>Tag1q =>L2Cmd =>Ipv4 =>Udp =>L3_1588);
    bins EthMacSec8VnTagTag1qL2CmdIpv6UdpL3_1588Trans = (Eth =>MacSec8 =>VnTag =>Tag1q =>L2Cmd =>Ipv6 =>Udp =>L3_1588);
    bins EthMacSec8VnTagTag1qL2CmdIpv6Ipv6ExtnDstnOption2UdpL3_1588Trans = (Eth =>MacSec8 =>VnTag =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Udp =>L3_1588);
    bins EthMacSec8VnTagTag1qL2CmdIpv6Ipv6ExtnFragmentUdpL3_1588Trans = (Eth =>MacSec8 =>VnTag =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Udp =>L3_1588);
    bins EthMacSec16Ipv4UdpL3_1588Trans = (Eth =>MacSec16 =>Ipv4 =>Udp =>L3_1588);
    bins EthMacSec16Ipv6UdpL3_1588Trans = (Eth =>MacSec16 =>Ipv6 =>Udp =>L3_1588);
    bins EthMacSec16Ipv6Ipv6ExtnDstnOption2UdpL3_1588Trans = (Eth =>MacSec16 =>Ipv6Ipv6ExtnDstnOption2 =>Udp =>L3_1588);
    bins EthMacSec16Ipv6Ipv6ExtnFragmentUdpL3_1588Trans = (Eth =>MacSec16 =>Ipv6Ipv6ExtnFragment =>Udp =>L3_1588);
    bins EthMacSec16L2CmdIpv4UdpL3_1588Trans = (Eth =>MacSec16 =>L2Cmd =>Ipv4 =>Udp =>L3_1588);
    bins EthMacSec16L2CmdIpv6UdpL3_1588Trans = (Eth =>MacSec16 =>L2Cmd =>Ipv6 =>Udp =>L3_1588);
    bins EthMacSec16L2CmdIpv6Ipv6ExtnDstnOption2UdpL3_1588Trans = (Eth =>MacSec16 =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Udp =>L3_1588);
    bins EthMacSec16L2CmdIpv6Ipv6ExtnFragmentUdpL3_1588Trans = (Eth =>MacSec16 =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Udp =>L3_1588);
    bins EthMacSec16Tag1qIpv4UdpL3_1588Trans = (Eth =>MacSec16 =>Tag1q =>Ipv4 =>Udp =>L3_1588);
    bins EthMacSec16Tag1qIpv6UdpL3_1588Trans = (Eth =>MacSec16 =>Tag1q =>Ipv6 =>Udp =>L3_1588);
    bins EthMacSec16Tag1qIpv6Ipv6ExtnDstnOption2UdpL3_1588Trans = (Eth =>MacSec16 =>Tag1q =>Ipv6Ipv6ExtnDstnOption2 =>Udp =>L3_1588);
    bins EthMacSec16Tag1qIpv6Ipv6ExtnFragmentUdpL3_1588Trans = (Eth =>MacSec16 =>Tag1q =>Ipv6Ipv6ExtnFragment =>Udp =>L3_1588);
    bins EthMacSec16Tag1qL2CmdIpv4UdpL3_1588Trans = (Eth =>MacSec16 =>Tag1q =>L2Cmd =>Ipv4 =>Udp =>L3_1588);
    bins EthMacSec16Tag1qL2CmdIpv6UdpL3_1588Trans = (Eth =>MacSec16 =>Tag1q =>L2Cmd =>Ipv6 =>Udp =>L3_1588);
    bins EthMacSec16Tag1qL2CmdIpv6Ipv6ExtnDstnOption2UdpL3_1588Trans = (Eth =>MacSec16 =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Udp =>L3_1588);
    bins EthMacSec16Tag1qL2CmdIpv6Ipv6ExtnFragmentUdpL3_1588Trans = (Eth =>MacSec16 =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Udp =>L3_1588);
    bins EthMacSec16VnTagTag1qIpv4UdpL3_1588Trans = (Eth =>MacSec16 =>VnTag =>Tag1q =>Ipv4 =>Udp =>L3_1588);
    bins EthMacSec16VnTagTag1qIpv6UdpL3_1588Trans = (Eth =>MacSec16 =>VnTag =>Tag1q =>Ipv6 =>Udp =>L3_1588);
    bins EthMacSec16VnTagTag1qIpv6Ipv6ExtnDstnOption2UdpL3_1588Trans = (Eth =>MacSec16 =>VnTag =>Tag1q =>Ipv6Ipv6ExtnDstnOption2 =>Udp =>L3_1588);
    bins EthMacSec16VnTagTag1qIpv6Ipv6ExtnFragmentUdpL3_1588Trans = (Eth =>MacSec16 =>VnTag =>Tag1q =>Ipv6Ipv6ExtnFragment =>Udp =>L3_1588);
    bins EthMacSec16VnTagTag1qL2CmdIpv4UdpL3_1588Trans = (Eth =>MacSec16 =>VnTag =>Tag1q =>L2Cmd =>Ipv4 =>Udp =>L3_1588);
    bins EthMacSec16VnTagTag1qL2CmdIpv6UdpL3_1588Trans = (Eth =>MacSec16 =>VnTag =>Tag1q =>L2Cmd =>Ipv6 =>Udp =>L3_1588);
    bins EthMacSec16VnTagTag1qL2CmdIpv6Ipv6ExtnDstnOption2UdpL3_1588Trans = (Eth =>MacSec16 =>VnTag =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnDstnOption2 =>Udp =>L3_1588);
    bins EthMacSec16VnTagTag1qL2CmdIpv6Ipv6ExtnFragmentUdpL3_1588Trans = (Eth =>MacSec16 =>VnTag =>Tag1q =>L2Cmd =>Ipv6Ipv6ExtnFragment =>Udp =>L3_1588);
    bins EthSapTrans = (Eth =>Sap);
    bins EthSnapTrans = (Eth =>Snap);
    bins EthTag1qSapTrans = (Eth =>Tag1q =>Sap);
    bins EthTag1qSnapTrans = (Eth =>Tag1q =>Snap);
    bins EthTag1qTag1qSapTrans = (Eth =>Tag1qTag1q =>Sap);
    bins EthTag1qTag1qSnapTrans = (Eth =>Tag1qTag1q =>Snap);
    bins EthStagSapTrans = (Eth =>Stag =>Sap);
    bins EthStagSnapTrans = (Eth =>Stag =>Snap);
    bins EthStagTag1qSapTrans = (Eth =>StagTag1q =>Sap);
    bins EthStagTag1qSnapTrans = (Eth =>StagTag1q =>Snap);
    bins EthVnTagTag1qSapTrans = (Eth =>VnTag =>Tag1q =>Sap);
    bins EthVnTagTag1qSnapTrans = (Eth =>VnTag =>Tag1q =>Snap);
    bins EthVnTagTag1qL2CmdSapTrans = (Eth =>VnTag =>Tag1q =>L2Cmd =>Sap);
    bins EthVnTagTag1qL2CmdSnapTrans = (Eth =>VnTag =>Tag1q =>L2Cmd =>Snap);
    bins EthMacSec8SapTrans = (Eth =>MacSec8 =>Sap);
    bins EthMacSec8SnapTrans = (Eth =>MacSec8 =>Snap);
    bins EthMacSec8L2CmdSapTrans = (Eth =>MacSec8 =>L2Cmd =>Sap);
    bins EthMacSec8L2CmdSnapTrans = (Eth =>MacSec8 =>L2Cmd =>Snap);
    bins EthMacSec8Tag1qSapTrans = (Eth =>MacSec8 =>Tag1q =>Sap);
    bins EthMacSec8Tag1qSnapTrans = (Eth =>MacSec8 =>Tag1q =>Snap);
    bins EthMacSec8Tag1qL2CmdSapTrans = (Eth =>MacSec8 =>Tag1q =>L2Cmd =>Sap);
    bins EthMacSec8Tag1qL2CmdSnapTrans = (Eth =>MacSec8 =>Tag1q =>L2Cmd =>Snap);
    bins EthMacSec8Tag1qTag1qSapTrans = (Eth =>MacSec8 =>Tag1qTag1q =>Sap);
    bins EthMacSec8Tag1qTag1qSnapTrans = (Eth =>MacSec8 =>Tag1qTag1q =>Snap);
    bins EthMacSec8Tag1qTag1qL2CmdSapTrans = (Eth =>MacSec8 =>Tag1qTag1q =>L2Cmd =>Sap);
    bins EthMacSec8Tag1qTag1qL2CmdSnapTrans = (Eth =>MacSec8 =>Tag1qTag1q =>L2Cmd =>Snap);
    bins EthMacSec8StagSapTrans = (Eth =>MacSec8 =>Stag =>Sap);
    bins EthMacSec8StagSnapTrans = (Eth =>MacSec8 =>Stag =>Snap);
    bins EthMacSec8StagL2CmdSapTrans = (Eth =>MacSec8 =>Stag =>L2Cmd =>Sap);
    bins EthMacSec8StagL2CmdSnapTrans = (Eth =>MacSec8 =>Stag =>L2Cmd =>Snap);
    bins EthMacSec8StagTag1qSapTrans = (Eth =>MacSec8 =>StagTag1q =>Sap);
    bins EthMacSec8StagTag1qSnapTrans = (Eth =>MacSec8 =>StagTag1q =>Snap);
    bins EthMacSec8StagTag1qL2CmdSapTrans = (Eth =>MacSec8 =>StagTag1q =>L2Cmd =>Sap);
    bins EthMacSec8StagTag1qL2CmdSnapTrans = (Eth =>MacSec8 =>StagTag1q =>L2Cmd =>Snap);
    bins EthMacSec8VnTagTag1qSapTrans = (Eth =>MacSec8 =>VnTag =>Tag1q =>Sap);
    bins EthMacSec8VnTagTag1qSnapTrans = (Eth =>MacSec8 =>VnTag =>Tag1q =>Snap);
    bins EthMacSec8VnTagTag1qL2CmdSapTrans = (Eth =>MacSec8 =>VnTag =>Tag1q =>L2Cmd =>Sap);
    bins EthMacSec8VnTagTag1qL2CmdSnapTrans = (Eth =>MacSec8 =>VnTag =>Tag1q =>L2Cmd =>Snap);
    bins EthMacSec16SapTrans = (Eth =>MacSec16 =>Sap);
    bins EthMacSec16SnapTrans = (Eth =>MacSec16 =>Snap);
    bins EthMacSec16L2CmdSapTrans = (Eth =>MacSec16 =>L2Cmd =>Sap);
    bins EthMacSec16L2CmdSnapTrans = (Eth =>MacSec16 =>L2Cmd =>Snap);
    bins EthMacSec16Tag1qSapTrans = (Eth =>MacSec16 =>Tag1q =>Sap);
    bins EthMacSec16Tag1qSnapTrans = (Eth =>MacSec16 =>Tag1q =>Snap);
    bins EthMacSec16Tag1qL2CmdSapTrans = (Eth =>MacSec16 =>Tag1q =>L2Cmd =>Sap);
    bins EthMacSec16Tag1qL2CmdSnapTrans = (Eth =>MacSec16 =>Tag1q =>L2Cmd =>Snap);
    bins EthMacSec16Tag1qTag1qSapTrans = (Eth =>MacSec16 =>Tag1qTag1q =>Sap);
    bins EthMacSec16Tag1qTag1qSnapTrans = (Eth =>MacSec16 =>Tag1qTag1q =>Snap);
    bins EthMacSec16Tag1qTag1qL2CmdSapTrans = (Eth =>MacSec16 =>Tag1qTag1q =>L2Cmd =>Sap);
    bins EthMacSec16Tag1qTag1qL2CmdSnapTrans = (Eth =>MacSec16 =>Tag1qTag1q =>L2Cmd =>Snap);
    bins EthMacSec16StagSapTrans = (Eth =>MacSec16 =>Stag =>Sap);
    bins EthMacSec16StagSnapTrans = (Eth =>MacSec16 =>Stag =>Snap);
    bins EthMacSec16StagL2CmdSapTrans = (Eth =>MacSec16 =>Stag =>L2Cmd =>Sap);
    bins EthMacSec16StagL2CmdSnapTrans = (Eth =>MacSec16 =>Stag =>L2Cmd =>Snap);
    bins EthMacSec16StagTag1qSapTrans = (Eth =>MacSec16 =>StagTag1q =>Sap);
    bins EthMacSec16StagTag1qSnapTrans = (Eth =>MacSec16 =>StagTag1q =>Snap);
    bins EthMacSec16StagTag1qL2CmdSapTrans = (Eth =>MacSec16 =>StagTag1q =>L2Cmd =>Sap);
    bins EthMacSec16StagTag1qL2CmdSnapTrans = (Eth =>MacSec16 =>StagTag1q =>L2Cmd =>Snap);
    bins EthMacSec16VnTagTag1qSapTrans = (Eth =>MacSec16 =>VnTag =>Tag1q =>Sap);
    bins EthMacSec16VnTagTag1qSnapTrans = (Eth =>MacSec16 =>VnTag =>Tag1q =>Snap);
    bins EthMacSec16VnTagTag1qL2CmdSapTrans = (Eth =>MacSec16 =>VnTag =>Tag1q =>L2Cmd =>Sap);
    bins EthMacSec16VnTagTag1qL2CmdSnapTrans = (Eth =>MacSec16 =>VnTag =>Tag1q =>L2Cmd =>Snap);
    bins EthItagInnerEthTrans = (Eth =>Itag =>InnerEth);
    bins EthItagL2SiaInnerEthTrans = (Eth =>Itag =>L2Sia =>InnerEth);
    bins EthBtagItagInnerEthTrans = (Eth =>BtagItag =>InnerEth);
    bins EthBtagItagL2SiaInnerEthTrans = (Eth =>BtagItag =>L2Sia =>InnerEth);
    bins EthSilTag1qItagInnerEthTrans = (Eth =>SilTag1q =>Itag =>InnerEth);
    bins EthSilTag1qItagL2SiaInnerEthTrans = (Eth =>SilTag1q =>Itag =>L2Sia =>InnerEth);
    bins EthSilTag1qBtagItagInnerEthTrans = (Eth =>SilTag1q =>BtagItag =>InnerEth);
    bins EthSilTag1qBtagItagL2SiaInnerEthTrans = (Eth =>SilTag1q =>BtagItag =>L2Sia =>InnerEth);
    bins EthFchItagInnerEthTrans = (Eth =>Fch =>Itag =>InnerEth);
    bins EthFchItagL2SiaInnerEthTrans = (Eth =>Fch =>Itag =>L2Sia =>InnerEth);
    bins EthFchBtagItagInnerEthTrans = (Eth =>Fch =>BtagItag =>InnerEth);
    bins EthFchBtagItagL2SiaInnerEthTrans = (Eth =>Fch =>BtagItag =>L2Sia =>InnerEth);
    bins EthMacSec8ItagInnerEthTrans = (Eth =>MacSec8 =>Itag =>InnerEth);
    bins EthMacSec8ItagL2SiaInnerEthTrans = (Eth =>MacSec8 =>Itag =>L2Sia =>InnerEth);
    bins EthMacSec8ItagL2CmdInnerEthTrans = (Eth =>MacSec8 =>Itag =>L2Cmd =>InnerEth);
    bins EthMacSec8ItagL2CmdL2SiaInnerEthTrans = (Eth =>MacSec8 =>Itag =>L2Cmd =>L2Sia =>InnerEth);
    bins EthMacSec8BtagItagInnerEthTrans = (Eth =>MacSec8 =>BtagItag =>InnerEth);
    bins EthMacSec8BtagItagL2SiaInnerEthTrans = (Eth =>MacSec8 =>BtagItag =>L2Sia =>InnerEth);
    bins EthMacSec8BtagItagL2CmdInnerEthTrans = (Eth =>MacSec8 =>BtagItag =>L2Cmd =>InnerEth);
    bins EthMacSec8BtagItagL2CmdL2SiaInnerEthTrans = (Eth =>MacSec8 =>BtagItag =>L2Cmd =>L2Sia =>InnerEth);
    bins EthMacSec8SilTag1qItagInnerEthTrans = (Eth =>MacSec8 =>SilTag1q =>Itag =>InnerEth);
    bins EthMacSec8SilTag1qItagL2SiaInnerEthTrans = (Eth =>MacSec8 =>SilTag1q =>Itag =>L2Sia =>InnerEth);
    bins EthMacSec8SilTag1qItagL2CmdInnerEthTrans = (Eth =>MacSec8 =>SilTag1q =>Itag =>L2Cmd =>InnerEth);
    bins EthMacSec8SilTag1qItagL2CmdL2SiaInnerEthTrans = (Eth =>MacSec8 =>SilTag1q =>Itag =>L2Cmd =>L2Sia =>InnerEth);
    bins EthMacSec8SilTag1qBtagItagInnerEthTrans = (Eth =>MacSec8 =>SilTag1q =>BtagItag =>InnerEth);
    bins EthMacSec8SilTag1qBtagItagL2SiaInnerEthTrans = (Eth =>MacSec8 =>SilTag1q =>BtagItag =>L2Sia =>InnerEth);
    bins EthMacSec8SilTag1qBtagItagL2CmdInnerEthTrans = (Eth =>MacSec8 =>SilTag1q =>BtagItag =>L2Cmd =>InnerEth);
    bins EthMacSec8SilTag1qBtagItagL2CmdL2SiaInnerEthTrans = (Eth =>MacSec8 =>SilTag1q =>BtagItag =>L2Cmd =>L2Sia =>InnerEth);
    bins EthMacSec16ItagInnerEthTrans = (Eth =>MacSec16 =>Itag =>InnerEth);
    bins EthMacSec16ItagL2SiaInnerEthTrans = (Eth =>MacSec16 =>Itag =>L2Sia =>InnerEth);
    bins EthMacSec16ItagL2CmdInnerEthTrans = (Eth =>MacSec16 =>Itag =>L2Cmd =>InnerEth);
    bins EthMacSec16ItagL2CmdL2SiaInnerEthTrans = (Eth =>MacSec16 =>Itag =>L2Cmd =>L2Sia =>InnerEth);
    bins EthMacSec16BtagItagInnerEthTrans = (Eth =>MacSec16 =>BtagItag =>InnerEth);
    bins EthMacSec16BtagItagL2SiaInnerEthTrans = (Eth =>MacSec16 =>BtagItag =>L2Sia =>InnerEth);
    bins EthMacSec16BtagItagL2CmdInnerEthTrans = (Eth =>MacSec16 =>BtagItag =>L2Cmd =>InnerEth);
    bins EthMacSec16BtagItagL2CmdL2SiaInnerEthTrans = (Eth =>MacSec16 =>BtagItag =>L2Cmd =>L2Sia =>InnerEth);
    bins EthMacSec16SilTag1qItagInnerEthTrans = (Eth =>MacSec16 =>SilTag1q =>Itag =>InnerEth);
    bins EthMacSec16SilTag1qItagL2SiaInnerEthTrans = (Eth =>MacSec16 =>SilTag1q =>Itag =>L2Sia =>InnerEth);
    bins EthMacSec16SilTag1qItagL2CmdInnerEthTrans = (Eth =>MacSec16 =>SilTag1q =>Itag =>L2Cmd =>InnerEth);
    bins EthMacSec16SilTag1qItagL2CmdL2SiaInnerEthTrans = (Eth =>MacSec16 =>SilTag1q =>Itag =>L2Cmd =>L2Sia =>InnerEth);
    bins EthMacSec16SilTag1qBtagItagInnerEthTrans = (Eth =>MacSec16 =>SilTag1q =>BtagItag =>InnerEth);
    bins EthMacSec16SilTag1qBtagItagL2SiaInnerEthTrans = (Eth =>MacSec16 =>SilTag1q =>BtagItag =>L2Sia =>InnerEth);
    bins EthMacSec16SilTag1qBtagItagL2CmdInnerEthTrans = (Eth =>MacSec16 =>SilTag1q =>BtagItag =>L2Cmd =>InnerEth);
    bins EthMacSec16SilTag1qBtagItagL2CmdL2SiaInnerEthTrans = (Eth =>MacSec16 =>SilTag1q =>BtagItag =>L2Cmd =>L2Sia =>InnerEth);
}
endgroup
