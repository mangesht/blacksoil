
function rawTask();
$display("Inside rawTask\n");
endfunction 
